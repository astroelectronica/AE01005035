.title KiCad schematic
.include "../models/C2012X7R2A104K125AA_p.mod"
.include "../models/C3216X5R1C106M160AA_p.mod"
.include "../models/C3216X7R2A105M160AA_p.mod"
.include "../models/MAX15007A.lib"
XU3 /VIN 0 C2012X7R2A104K125AA_p
V1 /VIN 0 {VSOURCE}
XU2 /VIN 0 C3216X7R2A105M160AA_p
XU4 /VOUT 0 C3216X5R1C106M160AA_p
R1 /VIN /EN {REN}
XU1 /VIN unconnected-_U1-Pad2_ /EN unconnected-_U1-Pad4_ 0 unconnected-_U1-Pad6_ unconnected-_U1-Pad7_ /VOUT MAX15007A
I1 /VOUT 0 {ILOAD}
XU5 /VOUT 0 C2012X7R2A104K125AA_p
.end
